LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-- ENCORDE ASCII CHE DA PRIORIT� A LF POI A CR ED INFINE SE ENTRAMBI 
--SONO A ZERO CONVERTE I DATI DI CAMPIONE E GLITCH NEI CARATTERI ASCII CORRISPONDENTI
ENTITY ENC_B_ASCII IS
PORT(
		CAMPIONE : IN STD_LOGIC;
		GLITCH : IN STD_LOGIC;
		LF : IN STD_LOGIC;
		CR : IN STD_LOGIC;
		CODE_ASCII : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0 )
		);
END ENC_B_ASCII;

ARCHITECTURE BEH OF ENC_B_ASCII IS


BEGIN 


PROCESS (CAMPIONE,GLITCH, LF, CR)
VARIABLE MUX_PILOT : STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN

--THIS SIGNAL TAKE FIRST CAMPIONE THEN GLITCH
MUX_PILOT := CAMPIONE & GLITCH;

IF (LF = '1') THEN 
-- TRASMETTO LF
CODE_ASCII <=  "00001010";
ELSIF (CR ='1') THEN 
--TRASMETTO CR
CODE_ASCII <=	"00001101";
ELSE 
C1 : CASE MUX_PILOT IS

	WHEN "00" => 
	--TRASMETTO 0
	CODE_ASCII <= "00110000";
	
	WHEN "10" =>
	--TRASMETTO 1
	CODE_ASCII <= "00110001";
	
	WHEN "11" =>
	--TRASMETTO X
	CODE_ASCII <= "01011000";
	
	WHEN "01" =>
	--TRASMETTO x
	CODE_ASCII <= "01111000";
	
	WHEN OTHERS => 
	--TRASMETTO E
   CODE_ASCII <= "01000101";
   
	END CASE C1;
	END IF;
	END PROCESS;
END BEH ;

library ieee;
use ieee.std_logic_1164.all;

ENTITY SAMPLER IS 
PORT (
EXT_IN : IN STD_LOGIC; 
CLK : IN STD_LOGIC ;
SAMPLE : IN STD_LOGIC;
nRESET: IN STD_LOGIC;
ASY_RISING : OUT STD_LOGIC;
ASY_FALLING : OUT STD_LOGIC;
ASY_GLITCH : BUFFER STD_LOGIC;
OUT_CAMPIONE : OUT STD_LOGIC; 
GLITCH : OUT STD_LOGIC
);
END SAMPLER;

ARCHITECTURE BEH OF SAMPLER IS
 
COMPONENT GLITCH_EVALUATOR IS 
PORT(
EXT_IN : IN STD_LOGIC; 
CLK : IN STD_LOGIC ;
SAMPLE : IN STD_LOGIC;
nRESET: IN STD_LOGIC;
ASY_RISING: BUFFER STD_LOGIC;
ASY_FALLING : BUFFER STD_LOGIC;
ASY_GLITCH : OUT STD_LOGIC
);
END COMPONENT;

COMPONENT D_FF 
   port
   (
      CLK : in std_logic;
      CLRN : in std_logic;
      ENA : in std_logic;      
      D : in std_logic;
      Q : out std_logic
   );
end COMPONENT ; 

BEGIN


GLITCH_EVALUATOR_0 :  GLITCH_EVALUATOR PORT MAP(
		EXT_IN => EXT_IN,
		CLK => CLK,
		SAMPLE => SAMPLE,
		nRESET => nRESET,
		ASY_RISING => ASY_RISING,
		ASY_FALLING => ASY_FALLING,
		ASY_GLITCH => ASY_GLITCH 
		);
		
CAMPIONAMENTO_IN : D_FF PORT MAP (
      CLK => CLK,
      CLRN => nRESET,
      ENA => SAMPLE,  
      D => EXT_IN,
      Q =>OUT_CAMPIONE
		);
		
CAMPIONAMENTO_GLITCH : D_FF PORT MAP (		
		CLK => CLK,
      CLRN => nRESET,
      ENA => SAMPLE,  
      D => ASY_GLITCH,
      Q => GLITCH
		);
		
END BEH ;
library ieee;
use ieee.std_logic_1164.all;

ENTITY GLITCH_EVALUATOR IS 
PORT(
EXT_IN : IN STD_LOGIC; 
CLK : IN STD_LOGIC ;
SAMPLE : IN STD_LOGIC;
nRESET: IN STD_LOGIC;
ASY_RISING: BUFFER STD_LOGIC;
ASY_FALLING : BUFFER STD_LOGIC;
ASY_GLITCH : OUT STD_LOGIC
);
END GLITCH_EVALUATOR;

ARCHITECTURE BEH OF GLITCH_EVALUATOR IS

component T_FF 
  port(
        CLK: in std_logic;
        nRESET: in std_logic;
        T: in std_logic;
        Q: buffer std_logic
      );
end component ;

COMPONENT POSITIVE_EDGE_DETECTOR 
PORT(
EXT_IN : IN STD_LOGIC; 
CLK : IN STD_LOGIC ;
ALTERNATE : IN STD_LOGIC;
nRESET: IN STD_LOGIC;
RISING : BUFFER STD_LOGIC
);
END COMPONENT;

COMPONENT NEGATIVE_EDGE_DETECTOR 
PORT(
EXT_IN : IN STD_LOGIC; 
CLK : IN STD_LOGIC ;
ALTERNATE : IN STD_LOGIC;
nRESET: IN STD_LOGIC;
FALLING : BUFFER STD_LOGIC
);
END COMPONENT;

SIGNAL ALTERNATE: STD_LOGIC;

BEGIN

TFF_ALTERNATE : T_FF  port map(
        CLK => CLK ,
        nRESET => nRESET,
        T => SAMPLE,
        Q => ALTERNATE
      );


POSITIVE_EDGE_DETECTOR_1 : POSITIVE_EDGE_DETECTOR PORT MAP (
			EXT_IN => EXT_IN,
			CLK => CLK ,
			ALTERNATE => ALTERNATE,
			nRESET => nRESET,
			RISING => ASY_RISING
);

NEGATIVE_EDGE_DETECTOR_1 : NEGATIVE_EDGE_DETECTOR PORT MAP(EXT_IN => EXT_IN,
			CLK => CLK ,
			ALTERNATE => ALTERNATE,
			nRESET => nRESET,
			FALLING => ASY_FALLING
);

ASY_GLITCH <= ASY_RISING AND ASY_FALLING ;

END BEH;
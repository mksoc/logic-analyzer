LIBRARY IEEE;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

entity TRIGGER IS
PORT ( 
			CLK,nRST    : IN  STD_LOGIC;
			COMP_VALUE  : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
			COND_VALUE  : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
			EN_MEM,EN_LOOK4TRIG  : IN  STD_LOGIC ;
			START_RQ    : OUT STD_LOGIC 
		);
		END TRIGGER ;
		
ARCHITECTURE BEH OF TRIGGER IS

COMPONENT D_FF 
   port
   (
      CLK : in std_logic;
      CLRN : in std_logic;
      ENA : in std_logic;      
      D : in std_logic;
      Q : out std_logic
   );
end  COMPONENT ;

COMPONENT COMPARATOR  
PORT (	ELM_1,ELM_2 : IN STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
         EN : IN STD_LOGIC ;
			EQUAL : OUT STD_LOGIC
			);
			END COMPONENT;
			
SIGNAL MEM_CONDITION : STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL TR_RES : STD_LOGIC;

BEGIN

REG: 
FOR I IN 7 DOWNTO 0 GENERATE
BEGIN
REGISTRO : D_FF PORT MAP (CLK,nRST,EN_MEM ,COND_VALUE(I),MEM_CONDITION(I));
END GENERATE REG ;

COM : COMPARATOR PORT MAP (MEM_CONDITION,COMP_VALUE,EN_LOOK4TRIG,START_RQ);


END BEH ;
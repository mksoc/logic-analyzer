LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FULL_SAMPLER IS 
PORT(
EXT_IN : IN STD_LOGIC_VECTOR ( 7 DOWNTO 0); 
CLK : IN STD_LOGIC ;
SAMPLE : IN STD_LOGIC;
nRESET: IN STD_LOGIC;

ASY_RISING : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0); 

ASY_FALLING : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0); 

ASY_GLITCH : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0);

OUT_CAMPIONE : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0); 
GLITCH : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0)
);
END FULL_SAMPLER;

ARCHITECTURE BEH OF FULL_SAMPLER IS 
COMPONENT SAMPLER 
PORT (
EXT_IN : IN STD_LOGIC; 
CLK : IN STD_LOGIC ;
SAMPLE : IN STD_LOGIC;
nRESET: IN STD_LOGIC;
ASY_RISING : OUT STD_LOGIC;
ASY_FALLING : OUT STD_LOGIC;
ASY_GLITCH : BUFFER STD_LOGIC;
OUT_CAMPIONE : OUT STD_LOGIC; 
GLITCH : OUT STD_LOGIC
);
END COMPONENT ;
BEGIN

GEN : FOR I IN 7 DOWNTO 0 GENERATE 
SAMPLER_I : SAMPLER PORT MAP 
(
EXT_IN  => EXT_IN(I),
CLK  => CLK,
SAMPLE  => SAMPLE,
nRESET  => nRESET,


ASY_RISING => ASY_RISING(I),
ASY_FALLING => ASY_FALLING(I),
ASY_GLITCH => ASY_GLITCH(I),

OUT_CAMPIONE => OUT_CAMPIONE(I),
GLITCH => GLITCH(I)
);
END GENERATE GEN;

END BEH;
LIBRARY IEEE;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPARATOR IS 
PORT (	ELM_1,ELM_2 : IN STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
			EN : IN STD_LOGIC ;
			EQUAL : OUT STD_LOGIC
			);
			END COMPARATOR ;
			
ARCHITECTURE BEH OF COMPARATOR IS

BEGIN

PROCESS (ELM_1,ELM_2,EN)
BEGIN
IF (ELM_1 = ELM_2) AND EN = '1' THEN 
EQUAL <= '1';
ELSE 
EQUAL <= '0';
END IF;
END PROCESS;
END BEH;